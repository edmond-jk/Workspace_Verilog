module aes_encipher_block (
	input wire			clk,
	input wire			reset_n,
	input wire			next,
	input wire [3:0]	round,
	input wire [127:0]	round_key,
	
	input wire [127:0]  in_block,
	output wire [127:0]	out_block,
	output wire			ready	
	);
	 
	 
endmodule